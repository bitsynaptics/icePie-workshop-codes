module led (
	output wire led_blue_n,
	output wire led_amber_n
);

assign led_blue_n = 1'b0;
assign led_amber_n = 1'b0;

endmodule